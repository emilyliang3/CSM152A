`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:28:25 03/19/2013 
// Design Name: 
// Module Name:    NERP_demo_top 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module NERP_demo_top(
	input wire clk,			//master clock = 100MHz
	input wire clr,			//right-most pushbutton for reset
	output wire [6:0] seg,	//7-segment display LEDs
	output wire [3:0] an,	//7-segment display anode enable
//	output wire dp,			//7-segment display decimal point
	output wire [2:0] red,	//red vga output - 3 bits
	output wire [2:0] green,//green vga output - 3 bits
	output wire [2:0] blue,	//blue vga output - 3 bits
	output wire hsync,		//horizontal sync out
	output wire vsync,			//vertical sync out
	input wire [9:0] X_POS,
	input wire [9:0] Y_POS,
	input wire [2:0] color,
	input wire tool_on,
	input wire size_sel
	);

// 7-segment clock interconnect
wire segclk;

// VGA display clock interconnect
wire dclk;

// disable the 7-segment decimal points
//assign dp = 1;

// generate 7-segment clock & display clock
clockdiv U1(
	.clk(clk),
	.clr(clr),
	.segclk(segclk),
	.dclk(dclk)
	);

// 7-segment display controller
segdisplay U2(
	.segclk(segclk),
	.clr(clr),
	.seg(seg),
	.an(an),
	.tool_on(tool_on),
	.size_sel(size_sel),
	.color(color)
	);

// VGA controller
//vga640x480 U3(
//    .clk(clk),
//	.dclk(dclk),
//	.clr(clr),
//	.hsync(hsync),
//	.vsync(vsync),
//	.red(red),
//	.green(green),
//	.blue(blue),
//	.X_POS(X_POS),
//	.Y_POS(Y_POS),
//	.color(color),
//	.tool_on(tool_on),
//	.size_sel(size_sel)
//	);

endmodule
