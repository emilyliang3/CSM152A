`timescale 1ns / 1ps

module property_ctrl(
    input clk,
    input [2:0] sw,
    output tool_active
    );
    
    // switch 0- when on, tool is active
    
    
    
endmodule
